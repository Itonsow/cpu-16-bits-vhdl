LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SignExtend IS
    PORT (
        A : IN STD_LOGIC_VECTOR (0 TO 4); --input
        X : OUT STD_LOGIC_VECTOR(0 TO 15));--dado extendido
END SignExtend;

ARCHITECTURE SE OF SignExtend IS
BEGIN
    X <= STD_LOGIC_VECTOR(RESIZE(SIGNED(A), X'LENGTH));
END;