LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Cpu IS
    GENERIC (DATA_SIZE : INTEGER := 16);--tamanho padrao do barramento
    PORT (
        CLOCK : IN STD_LOGIC; -clk
        INSTRUCTION_OUT_IFID : OUT STD_LOGIC_VECTOR(0 TO 15);--instrucao q ta no registrador if/id
        DEB_REGS_PC : OUT STD_LOGIC_VECTOR(0 TO 15);--valor pc
        DEB_CONTROL : OUT STD_LOGIC; --bit control
        DEB_ULA_IN_1 : OUT STD_LOGIC_VECTOR(0 TO 15); --A
        DEB_ULA_IN_2 : OUT STD_LOGIC_VECTOR(0 TO 15);--B
        DEB_OUT_ULA : OUT STD_LOGIC_VECTOR(0 TO 15);--resultado da ula

        DEB_SINAL_MUX_MEMWB : OUT STD_LOGIC; --bit memtoreg
        DEB_SINAL_REG_WRITE : OUT STD_LOGIC; --regwrite

        DEB_FILE_REG_1 : OUT STD_LOGIC_VECTOR(0 TO 15);--reg1
        DEB_FILE_REG_2 : OUT STD_LOGIC_VECTOR(0 TO 15);--reg2
        DEB_FILE_REG_3 : OUT STD_LOGIC_VECTOR(0 TO 15);--reg3
        DEB_FILE_REG_AUX : OUT STD_LOGIC --sinal pra escrita
    );
END Cpu;
ARCHITECTURE CPU OF Cpu IS

    -- ControlUnit
    COMPONENT ControlUnit
        PORT (
            WB : OUT STD_LOGIC_VECTOR(0 TO 1);--sinais wb
            MEM : OUT STD_LOGIC_VECTOR(0 TO 2);--sinais mem
            EX : OUT STD_LOGIC_VECTOR(0 TO 4);--sinais ex
            INSTRUCTION : IN STD_LOGIC_VECTOR(0 TO 15)--instru
        );
    END COMPONENT;

    -- AluControl
    COMPONENT AluControl
        PORT (
            ALU_OP : IN STD_LOGIC_VECTOR(0 TO 2);--bit vindo controlunit
            FUNCT : IN STD_LOGIC; --bit que vai ver c é add ou sub
            ULA_CODE : OUT STD_LOGIC_VECTOR(0 TO 1)
        );
    END COMPONENT;

    -- Mux_2para1_32b 
    COMPONENT Mux_2para1_32b
        PORT (
            CONTROL : IN STD_LOGIC;
            A : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
            B : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
            X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1)
        );
    END COMPONENT;

    -- Alu
    COMPONENT Alu
        PORT (
            A : IN STD_LOGIC_VECTOR(0 TO 15); --operando
            B : IN STD_LOGIC_VECTOR(0 TO 15);--operando
            ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1);--seleciona qual vai ser a instruçao
            ALU_OUT : OUT STD_LOGIC_VECTOR(0 TO 15);--resultado
            ZERO : OUT STD_LOGIC
        );
    END COMPONENT;

    -- Data Memory
    COMPONENT DataMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 15);--end
            CLOCK : IN STD_LOGIC;--clk
            MEM_WRITE : IN STD_LOGIC; --controle
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 15);
            MEM_READ : IN STD_LOGIC;
            READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    -- InstructionMemory
    COMPONENT InstructionMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 15);
            INSTRUCTION : OUT STD_LOGIC_VECTOR(0 TO 15) := "0000000000000000"
        );
    END COMPONENT;

    -- PCIncrement
    COMPONENT PCIncrement
        PORT (
            PC : IN STD_LOGIC_VECTOR (0 TO 15);
            X : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    -- Reg_Pipe_IFID
    COMPONENT Reg_Pipe_IFID
        PORT (
            CLOCK : IN STD_LOGIC;
            IN_PC_MAIS_4 : IN STD_LOGIC_VECTOR(0 TO 15);
            IN_INSTR_MEM : IN STD_LOGIC_VECTOR(0 TO 15);

            OUT_PC_MAIS_4 : OUT STD_LOGIC_VECTOR(0 TO 15);
            OUT_INSTR_MEM : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    -- Mux_2to1_5b
    COMPONENT Mux_2to1_5b
        PORT (
            CONTROL : IN STD_LOGIC;
            A : IN STD_LOGIC_VECTOR (0 TO 3);
            B : IN STD_LOGIC_VECTOR (0 TO 3);
            X : OUT STD_LOGIC_VECTOR (0 TO 3)
        );

    END COMPONENT;

    -- Reg_Pipe_IDEX
    COMPONENT Reg_Pipe_IDEX
        PORT (
            CLOCK : IN STD_LOGIC;
            IDEX_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            IDEX_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            IDEX_IN_EX : IN STD_LOGIC_VECTOR(0 TO 4);
            IDEX_IN_PC : IN STD_LOGIC_VECTOR(0 TO 15);
            IDEX_IN_READ1 : IN STD_LOGIC_VECTOR(0 TO 15);
            IDEX_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 15);
            IDEX_IN_IMED : IN STD_LOGIC_VECTOR(0 TO 15);
            IDEX_IN_RT : IN STD_LOGIC_VECTOR(0 TO 3);
            IDEX_IN_RD : IN STD_LOGIC_VECTOR(0 TO 3);

            IDEX_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            IDEX_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            IDEX_OUT_EX : OUT STD_LOGIC_VECTOR(0 TO 4);
            IDEX_OUT_PC : OUT STD_LOGIC_VECTOR(0 TO 15);
            IDEX_OUT_READ1 : OUT STD_LOGIC_VECTOR(0 TO 15);
            IDEX_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 15);
            IDEX_OUT_IMED : OUT STD_LOGIC_VECTOR(0 TO 15);
            IDEX_OUT_RT : OUT STD_LOGIC_VECTOR(0 TO 3);
            IDEX_OUT_RD : OUT STD_LOGIC_VECTOR(0 TO 3)
        );
    END COMPONENT;

    -- Reg_Pipe_EXMEM
    COMPONENT Reg_Pipe_EXMEM
        PORT (
            CLOCK : IN STD_LOGIC;
            EXMEM_IN_ZERO : IN STD_LOGIC;
            EXMEM_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_IN_RESULT_ADDER : IN STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 3);

            EXMEM_OUT_ZERO : OUT STD_LOGIC;
            EXMEM_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_OUT_RESULT_ADDER : OUT STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 15);
            EXMEM_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 3)
        );
    END COMPONENT;

    -- Reg_Pipe_MEMWB
    COMPONENT Reg_Pipe_MEMWB
        PORT (
            CLOCK : IN STD_LOGIC;
            MEMWB_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 15);
            MEMWB_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 3);
            MEMWB_IN_READ_DATA : IN STD_LOGIC_VECTOR(0 TO 15);

            MEMWB_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 15);
            MEMWB_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 3);
            MEMWB_OUT_READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    -- FileRegister
    COMPONENT FileRegister
        PORT (
            REGWRITE : IN STD_LOGIC;
            CLOCK : IN STD_LOGIC;
            READ_REGISTER_1 : IN STD_LOGIC_VECTOR(0 TO 3);
            READ_REGISTER_2 : IN STD_LOGIC_VECTOR(0 TO 3);
            WRITE_REGISTER : IN STD_LOGIC_VECTOR(0 TO 3);
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 15);

            READ_DATA_1 : OUT STD_LOGIC_VECTOR(0 TO 15);
            READ_DATA_2 : OUT STD_LOGIC_VECTOR(0 TO 15);

            DEB_FILE_REG_1 : OUT STD_LOGIC_VECTOR(0 TO 15);

            DEB_FILE_REG_2 : OUT STD_LOGIC_VECTOR(0 TO 15);
            DEB_FILE_REG_3 : OUT STD_LOGIC_VECTOR(0 TO 15);
            DEB_FILE_REG_AUX : OUT STD_LOGIC
        );
    END COMPONENT;

    -- ProgramCounter
    COMPONENT ProgramCounter
        PORT (
            CLOCK : IN STD_LOGIC;
            PC_INC : IN STD_LOGIC_VECTOR(0 TO 15);
            PC : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    -- SINAL EXTENDIDO
    COMPONENT SignExtend
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 4);
            X : OUT STD_LOGIC_VECTOR(0 TO 15)
        );
    END COMPONENT;

    --INSTRUCAO FETCH

    SIGNAL WIRE_OUT_PC_INC : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_OUT_PC : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_INST_MEM_IFID : STD_LOGIC_VECTOR(0 TO 15);
    
    --ESTAGIO DE DECODE
    SIGNAL WIRE_PC_INC_IFID_TO_IDEX : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_OUT_IFID_INSTRUCTION : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_READ_DATA1_IDEX : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_READ_DATA2_IDEX : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_SIGNAL_EXTEND_IDEX : STD_LOGIC_VECTOR(0 TO 15);

    --Control Unit
    SIGNAL WIRE_UC_IDEX_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_UC_IDEX_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_UC_IDEX_EX : STD_LOGIC_VECTOR(0 TO 4);

    --ESTAGIO DE EXECUCAO
    SIGNAL WIRE_IDEX_WB_EXMEM_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_IDEX_MEM_EXMEM_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_PC_INC_IDEX : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_IDEX_READ1_ALU_A : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_OUT_IDEX_READ2 : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_OUT_IDEX_IMED : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_IDEX_RT_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 3);
    SIGNAL WIRE_IDEX_RD_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 3);
    SIGNAL WIRE_OUT_IDEX_EX : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_MUX_ALU_B : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_MUX_REGDST_EXMEM : STD_LOGIC_VECTOR(0 TO 3);
    SIGNAL WIRE_ULA_CODE : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_ALU_RES_EXMEM : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_ZERO_EXMEM : STD_LOGIC;

    SIGNAL WIRE_OUT_EXMEM_ZERO : STD_LOGIC;
    SIGNAL WIRE_EXMEM_WB_MEMWB_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_OUT_EXMEM_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_OUT_EXMEM_ALU_RES : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_EXMEM_READ2_WRITE_DATA : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_EXMEM_REGDST_MEM_WB : STD_LOGIC_VECTOR(0 TO 3);

    SIGNAL WIRE_READ_DATA_MEMWB : STD_LOGIC_VECTOR(0 TO 15);

    --WRITE BACK ESTAGIO

    SIGNAL WIRE_OUT_MEMWB_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_MEMWB_ALU_RES : STD_LOGIC_VECTOR(0 TO 15);
    SIGNAL WIRE_MEMWB_REG_DST : STD_LOGIC_VECTOR(0 TO 3);
    SIGNAL WIRE_MEMWB_READ_DATA_MUX_WB : STD_LOGIC_VECTOR(0 TO 15);
    --
    SIGNAL WIRE_MUX_WB_WRITE_DATA : STD_LOGIC_VECTOR(0 TO 15);

BEGIN

    --FETCH

    INST_MEM : InstructionMemory PORT MAP(WIRE_OUT_PC, WIRE_INST_MEM_IFID);
    PC_INC : PCIncrement PORT MAP(WIRE_OUT_PC, WIRE_OUT_PC_INC);
    PC : ProgramCounter PORT MAP(CLOCK, WIRE_OUT_PC_INC, WIRE_OUT_PC);

    DEB_REGS_PC <= WIRE_OUT_PC_INC;
    --REG_PIPE IF/ID

    IFID : Reg_Pipe_IFID PORT MAP(CLOCK, WIRE_OUT_PC_INC, WIRE_INST_MEM_IFID, WIRE_PC_INC_IFID_TO_IDEX, WIRE_OUT_IFID_INSTRUCTION);

    INSTRUCTION_OUT_IFID <= WIRE_OUT_IFID_INSTRUCTION;

    --ESTAGIO DE DECODE 

    DEB_SINAL_REG_WRITE <= WIRE_OUT_MEMWB_WB(0);
    FILE_REG : FileRegister PORT MAP(
        WIRE_OUT_MEMWB_WB(0),
        CLOCK,
        WIRE_OUT_IFID_INSTRUCTION(3 TO 6),   -- RS: bits 3-6 (4 bits)
        WIRE_OUT_IFID_INSTRUCTION(7 TO 10),  -- RT: bits 7-10 (4 bits)
        WIRE_MEMWB_REG_DST,
        WIRE_MUX_WB_WRITE_DATA,
        WIRE_READ_DATA1_IDEX,
        WIRE_READ_DATA2_IDEX,

        DEB_FILE_REG_1,
        DEB_FILE_REG_2,
        DEB_FILE_REG_3,

        DEB_FILE_REG_AUX
    );
    SIGNAL_EXTEND : SignExtend PORT MAP(WIRE_OUT_IFID_INSTRUCTION(11 TO 15), WIRE_SIGNAL_EXTEND_IDEX);
    UC : ControlUnit PORT MAP(WIRE_UC_IDEX_WB, WIRE_UC_IDEX_MEM, WIRE_UC_IDEX_EX, WIRE_OUT_IFID_INSTRUCTION);

    --REG PIPE ID/EX
    IDEX : Reg_Pipe_IDEX PORT MAP(
        -- IN --
        CLOCK, WIRE_UC_IDEX_WB, WIRE_UC_IDEX_MEM, WIRE_UC_IDEX_EX, WIRE_PC_INC_IFID_TO_IDEX, WIRE_READ_DATA1_IDEX, WIRE_READ_DATA2_IDEX, WIRE_SIGNAL_EXTEND_IDEX, WIRE_OUT_IFID_INSTRUCTION(7 TO 10), WIRE_OUT_IFID_INSTRUCTION(11 TO 14),
        -- OUT --
        WIRE_IDEX_WB_EXMEM_WB, WIRE_IDEX_MEM_EXMEM_MEM, WIRE_OUT_IDEX_EX, WIRE_PC_INC_IDEX, WIRE_IDEX_READ1_ALU_A, WIRE_OUT_IDEX_READ2, WIRE_OUT_IDEX_IMED, WIRE_IDEX_RT_MUX_REGDST, WIRE_IDEX_RD_MUX_REGDST
    );
    --EXECUCAO

    MUX_ALU_B : Mux_2para1_32b PORT MAP(WIRE_OUT_IDEX_EX(4), WIRE_OUT_IDEX_READ2, WIRE_OUT_IDEX_IMED, WIRE_MUX_ALU_B);
    MUX_REGDST : Mux_2to1_5b PORT MAP(WIRE_OUT_IDEX_EX(0), WIRE_IDEX_RT_MUX_REGDST, WIRE_IDEX_RD_MUX_REGDST, WIRE_MUX_REGDST_EXMEM);
    ALU_CONTROL : AluControl PORT MAP(WIRE_OUT_IDEX_EX(1 TO 3), WIRE_OUT_IDEX_IMED(15), WIRE_ULA_CODE);
    MAIN_ALU : Alu PORT MAP(WIRE_IDEX_READ1_ALU_A, WIRE_MUX_ALU_B, WIRE_ULA_CODE, WIRE_ALU_RES_EXMEM, WIRE_ZERO_EXMEM);

    DEB_CONTROL <= WIRE_OUT_IDEX_EX(0);
    DEB_ULA_IN_1 <= WIRE_IDEX_READ1_ALU_A;
    DEB_ULA_IN_2 <= WIRE_MUX_ALU_B;
    DEB_OUT_ULA <= WIRE_ALU_RES_EXMEM;
    --REG_PIPE EX/MEM
    EXMEM : Reg_Pipe_EXMEM PORT MAP(
        -- IN --
        CLOCK,
        WIRE_ZERO_EXMEM,
        WIRE_IDEX_WB_EXMEM_WB,
        WIRE_IDEX_MEM_EXMEM_MEM,
        (OTHERS => '0'),  -- WIRE_ADDER_RES_EXMEM substituído por zeros (não usado)
        WIRE_ALU_RES_EXMEM,
        WIRE_OUT_IDEX_READ2,
        WIRE_MUX_REGDST_EXMEM,
        -- OUT --
        WIRE_OUT_EXMEM_ZERO,
        WIRE_EXMEM_WB_MEMWB_WB,
        WIRE_OUT_EXMEM_MEM,
        OPEN,  -- Resultado do adder não usado
        WIRE_OUT_EXMEM_ALU_RES,
        WIRE_EXMEM_READ2_WRITE_DATA,
        WIRE_EXMEM_REGDST_MEM_WB
    );

    DATA_MEMORY : DataMemory PORT MAP(WIRE_OUT_EXMEM_ALU_RES, CLOCK, WIRE_OUT_EXMEM_MEM(2), WIRE_EXMEM_READ2_WRITE_DATA, WIRE_OUT_EXMEM_MEM(1), WIRE_READ_DATA_MEMWB);

    --REG PIPE MEM/WB
    MEMWB : Reg_Pipe_MEMWB PORT MAP(
        -- IN --
        CLOCK,
        WIRE_EXMEM_WB_MEMWB_WB,
        WIRE_OUT_EXMEM_ALU_RES,
        WIRE_EXMEM_REGDST_MEM_WB,
        WIRE_READ_DATA_MEMWB,
        -- OUT --
        WIRE_OUT_MEMWB_WB,
        WIRE_MEMWB_ALU_RES,
        WIRE_MEMWB_REG_DST,
        WIRE_MEMWB_READ_DATA_MUX_WB
    );

    MUX_WB : Mux_2para1_32b PORT MAP(WIRE_OUT_MEMWB_WB(1), WIRE_MEMWB_READ_DATA_MUX_WB, WIRE_MEMWB_ALU_RES, WIRE_MUX_WB_WRITE_DATA);
    DEB_SINAL_MUX_MEMWB <= WIRE_OUT_MEMWB_WB(1);

END;