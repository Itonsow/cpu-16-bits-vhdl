LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ShiftLeft IS
    PORT (
        A : IN STD_LOGIC_VECTOR (0 TO 15);--DATA QUE VAI SER DESLOCADA
        X : OUT STD_LOGIC_VECTOR(0 TO 15)-- ONDE OS DADOS DESLOCADOS SAO ARMAZENADOS
    );
END ShiftLeft;

ARCHITECTURE SL OF ShiftLeft IS
BEGIN
    X <= A(1 TO 15) & "0"; -- Desloca 1 bit para esquerda (multiplica por 2)
END;