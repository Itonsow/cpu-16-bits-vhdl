LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PCincrement IS
    PORT (
        PC : IN STD_LOGIC_VECTOR (0 TO 15); --pc
        X : OUT STD_LOGIC_VECTOR(0 TO 15) := "0000000000000000");
END PCincrement;

ARCHITECTURE INC OF PCincrement IS
BEGIN
    X <= PC + "0000000000000010"; --pc+2
END;