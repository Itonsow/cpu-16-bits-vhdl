LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DataMemory IS
	PORT (
		ADDRESS : IN STD_LOGIC_VECTOR(0 TO 15);--endereco de acesso a memoria
		CLOCK : IN STD_LOGIC;
		MEM_WRITE : IN STD_LOGIC; --sinal de escrita
		WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 15); --oq vai ser escrito na memoria
		MEM_READ : IN STD_LOGIC;--sinal de leitura
		READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 15)); --lido da memoria

END DataMemory;

ARCHITECTURE MEM OF DataMemory IS
	TYPE MEM_TYPE IS ARRAY(0 TO 400) OF STD_LOGIC_VECTOR(0 TO 7);
	SIGNAL MEMORY : MEM_TYPE;
BEGIN
	PROCESS (CLOCK)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN
			IF (MEM_WRITE = '1') THEN --entra quando o sinal de escrita estiver ativo
				--Escreve 16 bits
				MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) <= WRITE_DATA(0 TO 7);
				MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1) <= WRITE_DATA(8 TO 15);
			END IF;

			IF (MEM_READ = '1') THEN
				-- Lê 16 bits (2 bytes)
				READ_DATA <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) &
					MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1);
			ELSE
				READ_DATA <= "ZZZZZZZZZZZZZZZZ";
			END IF;
		END IF;
	END PROCESS;
END;