LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

--operaçoes logicas

ENTITY Alu IS
	PORT (
		A : IN STD_LOGIC_VECTOR(0 TO 15);-- REGISTRADOR
		B : IN STD_LOGIC_VECTOR(0 TO 15); -- REGISTRADOR
		ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1); --CODIGO DA OPERACAO
		ALU_OUT : OUT STD_LOGIC_VECTOR(0 TO 15);-- ARMAZENAR O RESULTADO
		ZERO : OUT STD_LOGIC);
END Alu;

ARCHITECTURE ALU OF Alu IS
	SIGNAL AUX : STD_LOGIC_VECTOR(0 TO 15);
BEGIN
	PROCESS (A, B, ALU_CODE)
	BEGIN
		CASE ALU_CODE IS
			WHEN "00" => AUX <= A + B;--soma
			WHEN "01" => AUX <= A - B;--sub
			WHEN "10" => AUX <= A AND B; --and
			WHEN "11" => AUX <= A OR B;--or
			WHEN OTHERS => AUX <= "0000000000000000";
		END CASE;
		IF (AUX = "0000000000000000") THEN
			ZERO <= '1';
		ELSE
			ZERO <= '0';
		END IF;
		ALU_OUT <= AUX;
	END PROCESS;

END ALU;