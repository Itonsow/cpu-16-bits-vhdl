LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
--16
ENTITY Mux_2para1_32b IS
    GENERIC (DATA_SIZE : INTEGER := 16);
    PORT (
        CONTROL : IN STD_LOGIC;
        A : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
        B : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1); 
        X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1));
END Mux_2para1_32b;

ARCHITECTURE MUX OF Mux_2para1_32b IS
BEGIN
    X <= A WHEN (CONTROL = '0') ELSE B;
END;